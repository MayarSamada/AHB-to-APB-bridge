
module fsm ( Hclk, Hrstn, Hwrite, Hsel_APB, test_si, test_se, Haddr, Hwdata, 
        Prdata, Htrans, Hready_out, Penable, Pselx, Pwrite, test_so, Hrdata, 
        Pwdata, Paddr, Hresp );
  input [31:0] Haddr;
  input [31:0] Hwdata;
  input [31:0] Prdata;
  input [1:0] Htrans;
  output [31:0] Hrdata;
  output [31:0] Pwdata;
  output [31:0] Paddr;
  output [1:0] Hresp;
  input Hclk, Hrstn, Hwrite, Hsel_APB, test_si, test_se;
  output Hready_out, Penable, Pselx, Pwrite, test_so;
  wire   n46, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44,
         n45;
  wire   [2:0] current_state;
  wire   [2:0] next_state;
  assign Hresp[0] = 1'b0;
  assign Hresp[1] = 1'b0;

  DFFR_X1 current_state_reg_0_ ( .D(next_state[0]), .CK(Hclk), .RN(Hrstn), .Q(
        current_state[0]), .QN(n6) );
  DFFR_X1 current_state_reg_1_ ( .D(next_state[1]), .CK(Hclk), .RN(Hrstn), .Q(
        current_state[1]), .QN(n5) );
  DFFR_X1 current_state_reg_2_ ( .D(next_state[2]), .CK(Hclk), .RN(Hrstn), .Q(
        current_state[2]), .QN(n3) );
  INV_X1 U105 ( .A(n12), .ZN(n46) );
  INV_X1 U106 ( .A(n14), .ZN(n2) );
  INV_X1 U107 ( .A(n13), .ZN(n4) );
  INV_X1 U108 ( .A(n11), .ZN(n7) );
  NAND3_X1 U109 ( .A1(current_state[0]), .A2(n15), .A3(current_state[1]), .ZN(
        n8) );
  NAND3_X1 U110 ( .A1(n7), .A2(n6), .A3(Hwrite), .ZN(n10) );
  NAND2_X1 U111 ( .A1(Htrans[1]), .A2(Hsel_APB), .ZN(n11) );
  NAND2_X1 U112 ( .A1(n12), .A2(n13), .ZN(Pselx) );
  NAND2_X1 U113 ( .A1(current_state[2]), .A2(n5), .ZN(n12) );
  NAND2_X1 U114 ( .A1(current_state[0]), .A2(n5), .ZN(n13) );
  NAND2_X1 U115 ( .A1(n9), .A2(current_state[1]), .ZN(n14) );
  INV_X1 U116 ( .A(current_state[2]), .ZN(n15) );
  OR2_X1 U117 ( .A1(n9), .A2(Penable), .ZN(Hready_out) );
  OAI21_X1 U118 ( .B1(n5), .B2(n15), .A(n14), .ZN(Penable) );
  AND2_X1 U119 ( .A1(n3), .A2(n6), .ZN(n9) );
  AND2_X1 U120 ( .A1(Haddr[7]), .A2(n16), .ZN(Paddr[7]) );
  AND2_X1 U121 ( .A1(Haddr[8]), .A2(n16), .ZN(Paddr[8]) );
  AND2_X1 U122 ( .A1(Haddr[9]), .A2(n16), .ZN(Paddr[9]) );
  AND2_X1 U123 ( .A1(Haddr[1]), .A2(n21), .ZN(Paddr[1]) );
  AND2_X1 U124 ( .A1(Haddr[2]), .A2(n18), .ZN(Paddr[2]) );
  AND2_X1 U125 ( .A1(Haddr[3]), .A2(n17), .ZN(Paddr[3]) );
  AND2_X1 U126 ( .A1(Haddr[4]), .A2(n17), .ZN(Paddr[4]) );
  AND2_X1 U127 ( .A1(Haddr[5]), .A2(n17), .ZN(Paddr[5]) );
  AND2_X1 U128 ( .A1(Haddr[6]), .A2(n17), .ZN(Paddr[6]) );
  AND2_X1 U129 ( .A1(Haddr[10]), .A2(n23), .ZN(Paddr[10]) );
  AND2_X1 U130 ( .A1(Haddr[11]), .A2(n23), .ZN(Paddr[11]) );
  AND2_X1 U131 ( .A1(Haddr[12]), .A2(n23), .ZN(Paddr[12]) );
  AND2_X1 U132 ( .A1(Haddr[13]), .A2(n23), .ZN(Paddr[13]) );
  AND2_X1 U133 ( .A1(Haddr[14]), .A2(n22), .ZN(Paddr[14]) );
  AND2_X1 U134 ( .A1(Haddr[15]), .A2(n22), .ZN(Paddr[15]) );
  AND2_X1 U135 ( .A1(Haddr[16]), .A2(n22), .ZN(Paddr[16]) );
  AND2_X1 U136 ( .A1(Haddr[17]), .A2(n22), .ZN(Paddr[17]) );
  AND2_X1 U137 ( .A1(Haddr[18]), .A2(n21), .ZN(Paddr[18]) );
  AND2_X1 U138 ( .A1(Haddr[19]), .A2(n21), .ZN(Paddr[19]) );
  AND2_X1 U139 ( .A1(Haddr[20]), .A2(n21), .ZN(Paddr[20]) );
  AND2_X1 U140 ( .A1(Haddr[21]), .A2(n20), .ZN(Paddr[21]) );
  AND2_X1 U141 ( .A1(Haddr[22]), .A2(n20), .ZN(Paddr[22]) );
  AND2_X1 U142 ( .A1(Haddr[23]), .A2(n20), .ZN(Paddr[23]) );
  AND2_X1 U143 ( .A1(Haddr[24]), .A2(n20), .ZN(Paddr[24]) );
  AND2_X1 U144 ( .A1(Haddr[25]), .A2(n19), .ZN(Paddr[25]) );
  AND2_X1 U145 ( .A1(Haddr[26]), .A2(n19), .ZN(Paddr[26]) );
  AND2_X1 U146 ( .A1(Haddr[27]), .A2(n19), .ZN(Paddr[27]) );
  AND2_X1 U147 ( .A1(Haddr[28]), .A2(n19), .ZN(Paddr[28]) );
  AND2_X1 U148 ( .A1(Haddr[29]), .A2(n18), .ZN(Paddr[29]) );
  AND2_X1 U149 ( .A1(Haddr[30]), .A2(n18), .ZN(Paddr[30]) );
  AND2_X1 U150 ( .A1(Haddr[31]), .A2(n18), .ZN(Paddr[31]) );
  AND2_X1 U151 ( .A1(Hwdata[0]), .A2(n36), .ZN(Pwdata[0]) );
  AND2_X1 U152 ( .A1(Hwdata[1]), .A2(n38), .ZN(Pwdata[1]) );
  AND2_X1 U153 ( .A1(Hwdata[2]), .A2(n41), .ZN(Pwdata[2]) );
  AND2_X1 U154 ( .A1(Hwdata[3]), .A2(Pwrite), .ZN(Pwdata[3]) );
  AND2_X1 U155 ( .A1(Hwdata[4]), .A2(Pwrite), .ZN(Pwdata[4]) );
  AND2_X1 U156 ( .A1(Hwdata[5]), .A2(Pwrite), .ZN(Pwdata[5]) );
  AND2_X1 U157 ( .A1(Hwdata[6]), .A2(n43), .ZN(Pwdata[6]) );
  AND2_X1 U158 ( .A1(Hwdata[7]), .A2(n43), .ZN(Pwdata[7]) );
  AND2_X1 U159 ( .A1(Hwdata[8]), .A2(n43), .ZN(Pwdata[8]) );
  AND2_X1 U160 ( .A1(Hwdata[9]), .A2(n43), .ZN(Pwdata[9]) );
  AND2_X1 U161 ( .A1(Hwdata[10]), .A2(n36), .ZN(Pwdata[10]) );
  AND2_X1 U162 ( .A1(Hwdata[11]), .A2(n36), .ZN(Pwdata[11]) );
  AND2_X1 U163 ( .A1(Hwdata[12]), .A2(n36), .ZN(Pwdata[12]) );
  AND2_X1 U164 ( .A1(Hwdata[13]), .A2(n37), .ZN(Pwdata[13]) );
  AND2_X1 U165 ( .A1(Hwdata[14]), .A2(n37), .ZN(Pwdata[14]) );
  AND2_X1 U166 ( .A1(Hwdata[15]), .A2(n37), .ZN(Pwdata[15]) );
  AND2_X1 U167 ( .A1(Hwdata[16]), .A2(n37), .ZN(Pwdata[16]) );
  AND2_X1 U168 ( .A1(Hwdata[17]), .A2(n38), .ZN(Pwdata[17]) );
  AND2_X1 U169 ( .A1(Hwdata[18]), .A2(n38), .ZN(Pwdata[18]) );
  AND2_X1 U170 ( .A1(Hwdata[19]), .A2(n38), .ZN(Pwdata[19]) );
  AND2_X1 U171 ( .A1(Hwdata[20]), .A2(n39), .ZN(Pwdata[20]) );
  AND2_X1 U172 ( .A1(Hwdata[21]), .A2(n39), .ZN(Pwdata[21]) );
  AND2_X1 U173 ( .A1(Hwdata[22]), .A2(n39), .ZN(Pwdata[22]) );
  AND2_X1 U174 ( .A1(Hwdata[23]), .A2(n39), .ZN(Pwdata[23]) );
  AND2_X1 U175 ( .A1(Hwdata[24]), .A2(n40), .ZN(Pwdata[24]) );
  AND2_X1 U176 ( .A1(Hwdata[25]), .A2(n40), .ZN(Pwdata[25]) );
  AND2_X1 U177 ( .A1(Hwdata[26]), .A2(n40), .ZN(Pwdata[26]) );
  AND2_X1 U178 ( .A1(Hwdata[27]), .A2(n40), .ZN(Pwdata[27]) );
  AND2_X1 U179 ( .A1(Hwdata[28]), .A2(n41), .ZN(Pwdata[28]) );
  AND2_X1 U180 ( .A1(Hwdata[29]), .A2(n41), .ZN(Pwdata[29]) );
  AND2_X1 U181 ( .A1(Hwdata[30]), .A2(n41), .ZN(Pwdata[30]) );
  AND2_X1 U182 ( .A1(Hwdata[31]), .A2(Pwrite), .ZN(Pwdata[31]) );
  AND2_X1 U183 ( .A1(Prdata[0]), .A2(n26), .ZN(Hrdata[0]) );
  AND2_X1 U184 ( .A1(Prdata[1]), .A2(n28), .ZN(Hrdata[1]) );
  AND2_X1 U185 ( .A1(Prdata[2]), .A2(n31), .ZN(Hrdata[2]) );
  AND2_X1 U186 ( .A1(Prdata[3]), .A2(n32), .ZN(Hrdata[3]) );
  AND2_X1 U187 ( .A1(Prdata[4]), .A2(n32), .ZN(Hrdata[4]) );
  AND2_X1 U188 ( .A1(Prdata[5]), .A2(n32), .ZN(Hrdata[5]) );
  AND2_X1 U189 ( .A1(Prdata[6]), .A2(n33), .ZN(Hrdata[6]) );
  AND2_X1 U190 ( .A1(Prdata[7]), .A2(n33), .ZN(Hrdata[7]) );
  AND2_X1 U191 ( .A1(Prdata[8]), .A2(n33), .ZN(Hrdata[8]) );
  AND2_X1 U192 ( .A1(Prdata[9]), .A2(n33), .ZN(Hrdata[9]) );
  AND2_X1 U193 ( .A1(Prdata[10]), .A2(n26), .ZN(Hrdata[10]) );
  AND2_X1 U194 ( .A1(Prdata[11]), .A2(n26), .ZN(Hrdata[11]) );
  AND2_X1 U195 ( .A1(Prdata[12]), .A2(n26), .ZN(Hrdata[12]) );
  AND2_X1 U196 ( .A1(Prdata[13]), .A2(n27), .ZN(Hrdata[13]) );
  AND2_X1 U197 ( .A1(Prdata[14]), .A2(n27), .ZN(Hrdata[14]) );
  AND2_X1 U198 ( .A1(Prdata[15]), .A2(n27), .ZN(Hrdata[15]) );
  AND2_X1 U199 ( .A1(Prdata[16]), .A2(n27), .ZN(Hrdata[16]) );
  AND2_X1 U200 ( .A1(Prdata[17]), .A2(n28), .ZN(Hrdata[17]) );
  AND2_X1 U201 ( .A1(Prdata[18]), .A2(n28), .ZN(Hrdata[18]) );
  AND2_X1 U202 ( .A1(Prdata[19]), .A2(n28), .ZN(Hrdata[19]) );
  AND2_X1 U203 ( .A1(Prdata[20]), .A2(n29), .ZN(Hrdata[20]) );
  AND2_X1 U204 ( .A1(Prdata[21]), .A2(n29), .ZN(Hrdata[21]) );
  AND2_X1 U205 ( .A1(Prdata[22]), .A2(n29), .ZN(Hrdata[22]) );
  AND2_X1 U206 ( .A1(Prdata[23]), .A2(n29), .ZN(Hrdata[23]) );
  AND2_X1 U207 ( .A1(Prdata[24]), .A2(n30), .ZN(Hrdata[24]) );
  AND2_X1 U208 ( .A1(Prdata[25]), .A2(n30), .ZN(Hrdata[25]) );
  AND2_X1 U209 ( .A1(Prdata[26]), .A2(n30), .ZN(Hrdata[26]) );
  AND2_X1 U210 ( .A1(Prdata[27]), .A2(n30), .ZN(Hrdata[27]) );
  AND2_X1 U211 ( .A1(Prdata[28]), .A2(n31), .ZN(Hrdata[28]) );
  AND2_X1 U212 ( .A1(Prdata[29]), .A2(n31), .ZN(Hrdata[29]) );
  AND2_X1 U213 ( .A1(Prdata[30]), .A2(n31), .ZN(Hrdata[30]) );
  AND2_X1 U214 ( .A1(Prdata[31]), .A2(n32), .ZN(Hrdata[31]) );
  AND2_X1 U215 ( .A1(Haddr[0]), .A2(n4), .ZN(Paddr[0]) );
  OAI22_X1 U216 ( .A1(n16), .A2(n11), .B1(n6), .B2(n15), .ZN(next_state[0]) );
  OAI21_X1 U217 ( .B1(current_state[1]), .B2(n15), .A(n8), .ZN(next_state[2])
         );
  OAI21_X1 U218 ( .B1(current_state[1]), .B2(n9), .A(n10), .ZN(next_state[1])
         );
  INV_X1 U219 ( .A(n25), .ZN(n16) );
  INV_X1 U220 ( .A(n25), .ZN(n17) );
  INV_X1 U221 ( .A(n25), .ZN(n18) );
  INV_X1 U222 ( .A(n24), .ZN(n19) );
  INV_X1 U223 ( .A(n24), .ZN(n20) );
  INV_X1 U224 ( .A(n24), .ZN(n21) );
  INV_X1 U225 ( .A(n24), .ZN(n22) );
  INV_X1 U226 ( .A(n25), .ZN(n23) );
  INV_X1 U227 ( .A(n4), .ZN(n24) );
  INV_X1 U228 ( .A(n4), .ZN(n25) );
  INV_X1 U229 ( .A(n14), .ZN(n26) );
  INV_X1 U230 ( .A(n14), .ZN(n27) );
  INV_X1 U231 ( .A(n35), .ZN(n28) );
  INV_X1 U232 ( .A(n35), .ZN(n29) );
  INV_X1 U233 ( .A(n35), .ZN(n30) );
  INV_X1 U234 ( .A(n34), .ZN(n31) );
  INV_X1 U235 ( .A(n34), .ZN(n32) );
  INV_X1 U236 ( .A(n34), .ZN(n33) );
  INV_X1 U237 ( .A(n2), .ZN(n34) );
  INV_X1 U238 ( .A(n2), .ZN(n35) );
  INV_X1 U239 ( .A(n45), .ZN(n36) );
  INV_X1 U240 ( .A(n45), .ZN(n37) );
  INV_X1 U241 ( .A(n45), .ZN(n38) );
  INV_X1 U242 ( .A(n44), .ZN(n39) );
  INV_X1 U243 ( .A(n44), .ZN(n40) );
  INV_X1 U244 ( .A(n44), .ZN(n41) );
  INV_X1 U245 ( .A(n12), .ZN(Pwrite) );
  INV_X1 U246 ( .A(n12), .ZN(n43) );
  INV_X1 U247 ( .A(n46), .ZN(n44) );
  INV_X1 U248 ( .A(n46), .ZN(n45) );
endmodule

